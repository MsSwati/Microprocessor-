*OPAMP GENERATOR 
X1 1 0 5 6 2 UA741
.LIB UA741.LIB
VCC 5 0 DC 15V
VEE 0 6 DC 15V
Vin 1 0 ac 100v
R 2 0 0.001K 
.ac dec 100HZ 100HZ 1MegHz
.probe
.end